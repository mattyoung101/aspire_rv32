`default_nettype none

// This module decodes and expands RV32C compressed instructions.
