// This module implements Aspire's register file for FPGA.
// The implementation would be different for an ASIC.
