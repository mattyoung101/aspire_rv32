// This module implements Aspire's memory for an FPGA. Tries to make use of BRAM where possible.
