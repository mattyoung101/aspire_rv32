// The prefetcher communicates with the Winbond SPI flash to copy the program into the FPGA BRAM.
// Not required for simulation.
// For an ASIC tapeout, this module may require modification depending on how the SRAM cells
// are implemented.
