`default_nettype none

// This module implements Aspire's ALU.
