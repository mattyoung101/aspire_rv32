// Decoder for RV32I_Zmmul_Zicsr
