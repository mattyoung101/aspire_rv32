// Decoder for RV32IC_Zmmul_Zicsr
